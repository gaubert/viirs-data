netcdf GOME_NETCDF4 {

group: StatusData {
   
    group: SatelliteStatus {
	      :x_velocity=1418.549 ; // m/s
	      :y_velocity=848.027  ; // m/s
	      :z_velocity=7355.376 ; // m/s
	      :z_position=4865.973 ; // m
	      :x_position=-3742784.424 ; // m
	      :y_position=6152574.206 ; // m
		  :semi_major_axis=7204683346; // mm
		  :inclination=98.715; // deg
		  :eccentricity=0.00113;
		  :perigee_argument=67.634 ;//deg
		  :right_ascension=25.5 ;// deg
		  :mean_anomaly=292.525 ;// deg
		  :earth_sun_distance_ratio=6 ;//deg
		  :location_tolerance_radial=0 ;//m
		  :location_tolerance_crosstrack=0 ;//m
		  :location_tolerance_alongtrack=0; //m
		  :yaw_error=0; //deg
		  :roll_error=0; //deg
		  :pitch_error=0; //deg
		  :subsat_latitude_start=-81.314; //deg
		  :subsat_longitude_start=-164.53; //deg
		  :subsat_latitude_end=-76.716; //deg
		  :subsat_longitude_end=141.858; //deg	
    }

    group: InstrumentStatus {
	      :instrument_id="gome";
		  :instrument_model=1;
		  :processing_level="level 1b";
		  :spacecraft_id="m02";
		  :sensing_start="2010/11/24 14:38:58.000";
		  :sensing_end="2010/11/24 14:41:58.000";
		  :sensing_start_theoretical="2010/11/24 13:54:00.000";
		  :sensing_end_theoretical="2010/11/24 15:33:00.000";
    }

    group: ProcessingStatus {
	:MyGroup="1";
    }

}

group: MetaData { // Aux info

}

group: ScienceData {

	group: Product {

	dimensions:
		mdrs                     = 30; // Nb of MDRs in this file
		nb_pixels                = UNLIMITED;
		time                     = 1;
		pixels_4_itime_1.5       = 4;
		pixels_4_itime_6         = 1;
		pixels_4_itime_0.1875    = 32;
		pixels_4_itime_0.0234375 = 256;
		corners                  = 4; // nb of corners
		// number of elements per bands
		rec_band_1A              = 659;  // seems to be fix for all band_1A recs if not they should be defined locally in each group
		rec_band_1B              = 365;  // same
		rec_band_2A              = 71;   // same
		rec_band_2B              = 953;  // same
		rec_band_3               = 1024; // same
		rec_band_4               = 1024; // same
		rec_band_5               = 15;   // same
		rec_band_6               = 15;   // same
		rec_band_shortPS         = 20;   // same
		rec_band_shortPP         = 20;   // same
		nb_itimes                = 6;    // max number of integration times
		unknown_dim = 3; // do not know why it is always 3

	variables:
		// in this case itimes will always be the max possible 6 and the number of pixels will be the max for all MDRs. The number of pixels used will determine which integration time had been used
		// the maximum integration time used for all MDRs in this file is for example 0.1875 which means that we need to have nb_pixels = 32 
		// Fill values are also going to be used a lot and the file size will be a little bit inflated but compression should be good.
		int start_time(mdrs,time) ;
			start_time:long_name = "reference time of a MDR" ;
			start_time:units     = "UTC time in epoch time: seconds since 1971 (epoc time)" ;

		int end_time(mdrs,time) ;
			end_time:long_name = "reference time of a MDR" ;
			end_time:units     = "UTC time in epoch time: seconds since 1971 (epoc time): seconds since 1971 (epoc time)" ;

		float itimes(mdrs, nb_itimes); // integration times
			itimes:long_name = "integration times";
			itimes:units     = "seconds" ;
			itimes:_FillValue = -999 ;
			itimes:valid_min = -127b ;
			itimes:valid_max = 127b ;

		float scanner_angle(mdrs, nb_itimes, pixels_4_itime_0.1875); // take the max of nb pixels for all possible integration times, need to use invalid values for not existing values
			scanner_angle:long_name  = "scanner angle";
			scanner_angle:units      = "degrees" ;
			scanner_angle:_FillValue = -999 ; 
			scanner_angle:valid_min  = -180 ; // QC values (example, not the right values)
			scanner_angle:valid_max  = 180  ; // QC values (example, not the right values)
	  
		float corners(mdrs, nb_itimes, corners, pixels_4_itime_0.1875); // take the max of nb pixels for all possible integration times, need to use invalid values for not existing values
			corners:long_name   = "pixel corners";
			corners:units       = "degrees";
			corners:_FillValue  = -999;
			corners:valid_min   = -180; // QC values (example, not the right values) 
			corners:valid_max   = 180; // QC values (example, not the right values) 

		float centers(mdrs, nb_itimes, pixels_4_itime_0.1875); // take the max of nb pixels for all possible integration times, need to use invalid values for not existing values (here it is 32 values)
			corners:long_name   = "pixel centre";
			corners:units       = "degrees";
			corners:_FillValue  = -999;
			corners:valid_min   = -180; // QC values (example, not the right values) 
			corners:valid_max   = 180; // QC values (example, not the right values) 

		float solar_zenith(mdrs, nb_itimes, unknown_dim, pixels_4_itime_0.1875); // same take the max possible number of pixels for all possible integration times (here 32 values)
			solar_zenith:long_name  = "solar zenith";
			solar_zenith:units      = "degrees";
			solar_zenith:_FillValue = -999;
			solar_zenith:valid_min  = -180; // QC values (example, not the right values) 
			solar_zenith:valid_max  = 180; // QC values (example, not the right values) 

		float wavelength_1A(mdrs, rec_band_1A);
			wavelength_1A:long_name  = "wavelength values for band 1A";
			wavelength_1A:units      = "nm";  
			wavelength_1A:_FillValue = -9999; // TBD
			wavelength_1A:valid_min  = 0; // TBD 
			wavelength_1A:valid_max  = 0; // TBD 

		float band_1A(mdrs, pixels_4_itime_0.1875, rec_band_1A); //a band is nb of pixels * nb of measures in a record
			band_1A:long_name  = "measures for band 1A";
			band_1A:units      = "BU";  // TBD
			band_1A:_FillValue = -9999; // TBD
			band_1A:valid_min  = 0; // TBD 
			band_1A:valid_max  = 0; // TBD 

		float wavelength_1B(mdrs, rec_band_1B);
			wavelength_1B:long_name  = "wavelength values for band 1B";
			wavelength_1B:units      = "nm";  
			wavelength_1B:_FillValue = -9999; // TBD
			wavelength_1B:valid_min  = 0; // TBD 
			wavelength_1A:valid_max  = 0; // TBD 

		float band_1B(mdrs, pixels_4_itime_0.1875,rec_band_1B); //a band is nb of pixels * nb of measures in a record
			band_1B:long_name  = "measures for band 1B";
			band_1B:units      = "BU";  // TBD
			band_1B:_FillValue = -9999; // TBD
			band_1B:valid_min  = 0; // TBD 
			band_1B:valid_max  = 0; // TBD 

		// Add the other bands
	  } // group Product
  } // Science Data

// global attributes:
 :Conventions = "CF-1.0" ;
 :title = "GOME ..." ;
 :DSD_entry_id = "" ;
 :references = "N/A" ;
 :institution = "EUMETSAT:copyright 2011 EUMETSAT" ;
 :contact = "Eumetsat help desk at http://www.eumetsat.int" ;
 :netcdf_version_id = "netcdf library version 4.1.1 of Dec  2 2010 14:09:08" ;
 :creation_date = "2011-04-29" ;
 :product_version = "0.2" ;
}
