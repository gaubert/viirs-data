netcdf GOME_NETCDF4 {
types:
     compound f_range_t {
	     float start ;
	     float end ;
};

group: StatusData {

   // Remarques using attributes, we loose the unit
   // Metadata group is confusing because the netcdf header is already called metadata and the rest is also metadata data
   
   :spacecraft_id="m02";

   // Do not know where to put this information
   // Where to put that ?
  :duration_of_product_in_ms=180000; //ms
  :milliseconds_of_data_present=180000; //ms
  :milliseconds_of_data_missing=0; //ms

    group: SatelliteStatus {
		  :state_vector_time="2010-11-24T13:23:08.000Z";// ISO 8601 TIME
		  :orbit_start      =21266;
		  :orbit_stop       =21267;

	 variables:
	    float x_velocity;
	          x_velocity:units       = "m/s";
	          x_velocity:long_name   = "velocity on the x axis";
	    float y_velocity;
	          y_velocity:units       = "m/s";
	          y_velocity:long_name   = "velocity on the y axis";
	    float z_velocity;
	          z_velocity:units       = "m/s";
	          z_velocity:long_name   = "velocity on the z axis";
	    float x_position;
	          x_position:units       = "m";
	          x_position:long_name   = "satellite position on the x axis";
	    float y_position;
	          y_position:units       = "m";
	          y_position:long_name   = "satellite position on the y axis";
	    float z_position;
	          z_position:units       = "m";
	          z_position:long_name   = "satellite position on the z axis";
	    int   semi_major_axis;
	          semi_major_axis:units       = "mm";
	          semi_major_axis:long_name   = "semi major axis";
	    float inclination;
	          inclination:units       = "degrees";
	          inclination:long_name   = "satellite inclination";
	    float eccentricity;
	          eccentricity:units       = "degrees";
	          eccentricity:long_name   = "satellite eccentricity";
	    float perigee_argument;
	          perigee_argument:units       = "degrees";
	          perigee_argument:long_name   = "perigee argument";
	    float right_ascension;
	          right_ascension:units       = "degrees";
	          right_ascension:long_name   = "right ascension";
	    float mean_anomaly;
	          mean_anomaly:units       = "degrees";
	          mean_anomaly:long_name   = "mean anomaly";
        float earth_sun_distance_ratio;
	          earth_sun_distance_ratio:units            = "degrees";
			  earth_sun_distance_ratio:long_name        = "earth sun distance ratio";
	    float location_tolerance_radial;
	          location_tolerance_radial:units           = "degrees";
			  location_tolerance_radial:long_name       = "location tolerance radial";
        float location_tolerance_crosstrack;
	          location_tolerance_crosstrack:units       = "m";
			  location_tolerance_crosstrack:long_name   = "location tolerance crosstrack";
        float location_tolerance_alongtrack;
	          location_tolerance_alongtrack:units       = "m";
			  location_tolerance_alongtrack:long_name   = "location tolerance along track";
        float yaw_error;
	          yaw_error:units                           = "degrees";
			  yaw_error:long_name                       = "yaw error";
        float roll_error;
	          roll_error:units                          = "degrees";
			  roll_error:long_name                      = "roll error";
        float pitch_error;
	          pitch_error:units                         = "degrees";
			  pitch_error:long_name                     = "roll error";
        f_range_t subsat_latitude;
	          subsat_latitude:units                     = "degrees";
			  subsat_latitude:long_name                 = "subsatellite latitude start and end";
        f_range_t subsat_longitude;
	          subsat_longitude:units                    = "degrees";
			  subsat_longitude:long_name                = "subsatellite longitude start and end";
	           
	 data:
	     x_velocity                    = 1418.549;
	     y_velocity                    = 848.027;
	     z_velocity                    = 7355.376;
	     x_position                    = 4865.973;
	     y_position                    = 6152574.206;
	     z_position                    = -3742784.424;
		 semi_major_axis               = 7204683346;
		 perigee_argument              = 67.634;
		 inclination                   = 98.715;
		 eccentricity                  = 0.00113;
		 right_ascension               = 25.5;
		 mean_anomaly                  = 292.525;
		 location_tolerance_crosstrack =0;
		 location_tolerance_alongtrack =0;
		 yaw_error                     =0; 
		 roll_error                    =0; 
		 pitch_error                   =0;
		 subsat_latitude               = {-81.314, -76.716};
		 subsat_longitude              = {-164.53, 141.858};


    }

    group: InstrumentStatus {
	      :instrument_id="gome";
		  :instrument_model=1;
		  :processing_level="level 1b";
		  :sensing_start="2010-11-24T14:38:58.000Z"; //ISO TIME
		  :sensing_end="2010-11-24T14:41:58.000Z"; //ISO TIME
		  :sensing_start_theoretical="2010-11-24T13:54:00.000Z";
		  :sensing_end_theoretical="2010-11-24T15:33:00.000Z";
		  :leap_second=0;
		  :leap_second_utc="2013-06-19T10:34:30.296Z";

           
		  :n_scans=30; 
		  :n_valid_with_miss_dp=0; 
		  :n_miss_dp=0;
		  :n_missing_scans=0; 
		  :n_nn_detector_temp_1=0 ;
		  :n_nn_detector_temp_2=0 ;
          :n_nn_detector_temp_3=0 ;
    	  :n_nn_detector_temp_4=0 ;
		  :n_nn_detector_temp_5=0 ;
		  :n_nn_detector_temp_6=0 ;
		  :n_nn_pdp_temp=0 ;
		  :n_nn_rad_temp=0 ;
	  	  :n_nn_wls_u=0 ;
			:n_nn_wls_i=0 ;
			:n_nn_sls_u=0 ;
			:n_nn_sls_i=0 ;
			:n_inv_utc=0 ;
			:n_nadir_scan=30 ;
			:n_nth_pole_scan=0 ;
			:n_sth_pole_scan=0 ;
			:n_other_scan=0 ;
			:n_nadir_static=0 ;
			:n_other_static=0 ;
			:n_dark=0 ;
			:n_led=0 ;
			:n_wls=0 ;
			:n_sls=0 ;
			:n_sls_diff=0 ;
			:n_sun=0 ;
			:n_moon=0 ;
			:n_idle=0 ;
			:n_test=0 ;
			:n_dump=0 ;
			:n_invalid=0 ;
			:n_min_intensity_1=0 ;
			:n_min_intensity_2=0 ;
			:n_min_intensity_3=0 ;
			:n_min_intensity_4=0 ;
			:n_min_intensity_5=0 ;
			:n_min_intensity_6=0 ;
			:n_min_intensity_7=0 ;
			:n_min_intensity_8=0 ;
			:n_saturated_1=0 ;
			:n_saturated_2=0 ;
			:n_saturated_3=0 ;
			:n_saturated_4=0 ;
			:n_saturated_5=0 ;
			:n_saturated_6=0 ;
			:n_saturated_7=0 ;
			:n_saturated_8=0 ;
			:n_hot_1=0;
			:n_hot_2=0; 
			:n_hot_3=0; 
			:n_hot_4=0; 
			:n_hot_5=0; 
			:n_hot_6=0; 
			:n_hot_7=0; 
			:n_hot_8=0; 
			:n_saa=0; 
			:n_sunglint=0; 
			:n_rainbow=0; 
			:n_mode_geolocation=0; 
			:n_miss_stokes_1=11; 
			:n_miss_stokes_2=1; 
			:n_miss_stokes_3=0; 
			:n_miss_stokes_4=0; 
			:n_miss_stokes_5=0; 
			:n_miss_stokes_6=0; 
			:n_miss_stokes_7=0; 
			:n_miss_stokes_8=0; 
			:n_miss_stokes_9=0; 
			:n_miss_stokes_10=0; 
			:n_miss_stokes_11=0; 
			:n_miss_stokes_12=0; 
			:n_miss_stokes_13=0; 
			:n_miss_stokes_14=0; 
			:n_miss_stokes_15=0; 
			:n_bad_stokes_1=0; 
			:n_bad_stokes_2=0; 
			:n_bad_stokes_3=0; 
			:n_bad_stokes_4=0; 
			:n_bad_stokes_5=0; 
			:n_bad_stokes_6=0; 
			:n_bad_stokes_7=0; 
			:n_bad_stokes_8=0; 
			:n_bad_stokes_9=0; 
			:n_bad_stokes_1=0; 
			:n_bad_stokes_1=0; 
			:n_bad_stokes_1=0; 
			:n_bad_stokes_1=0; 
			:n_bad_stokes_14=0; 
			:n_bad_stokes_15=0; 
			:n_cloud=17; 
			:processing_indicator="xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx";
    }

    group: ProcessingStatus {
	      :processing_centre="cgs1";
		  :processor_major_version=4; 
		  :processor_minor_version=5; 
		  :format_major_version=11; 
		  :format_minor_version=0; 
		  :processing_time_start="2010-11-24T16:10:22.000Z"; // ISO 8601 TIME
		  :processing_time_end="2010-11-24T16:10:39.000Z"; // ISO 8601 TIME
		  :processing_mode="n"; 
    }
}

group: MetaData { // Would prefer to call it AuxiliaryData as MetaData is confusing

   :elevation="GOME_STA_xx_xxx_20070504000000Z_xxxxxxxxxxxxxxZ_20070503000103Z_xxxx_xxxxxxxxxx";

   :intialisation="GOME_INS_xx_M02_20100806000000Z_20251231235959Z_20100806000124Z_xxxx_FM3x440xxx";

   :keydata="GOME_CAL_xx_M02_20091105000000Z_xxxxxxxxxxxxxxZ_20091105000108Z_xxxx_FM3x440xxx";

 group: Channel {

	 dimensions:
		  chan_nb = 6;

	 variables:
		  f_range_t wave_length_range(chan_nb);
			 wave_length_range:long_name = "Wave length range for each channel" ;
			 wave_length_range:units     = "nm";

		  f_range_t valid_pixel_range(chan_nb);
			 valid_pixel_range:long_name = "pixel number for each channel" ;
			 valid_pixel_range:units     = "pixel position";
	
	  

	  data:
		 wave_length_range = { 239, 313.77}, { 309.45, 401.77}, { 395.35, 604.35}, { 592.56, 791}, {290,870}, {290,870};
		 valid_pixel_range = { 272, 942}, {151, 932}, {18, 1009}, {35, 989}, {750, 999}, {749, 1000};
}

group: Band1B {

	 dimensions:
		  chan_nb = 10;
		  band_nb = 10;

	 variables:

	      int chan_nb(chan_nb);
	         chan_nb:long_name = "Channel number";
		  int band_nb(band_nb);
	         band_nb:long_name = "Band number";

          int start_pixel(chan_nb);
	         start_pixel:long_name = "Start pixels of the different bands";

          int number_of_pixels(chan_nb);
	         number_of_pixels:long_name = "Number of pixels of the different bands";


		  f_range_t lambda_range(chan_nb);
			 lambda_range:long_name = "Wave length range for each channel" ;
			 lambda_range:units     = "nm";
 }

 // group 1b-steps
 // group 1b-pmdbandref
 // add viadr =>  time is used add the variable it qualifies and the time for which it is valid. Add attributes to qualify it 

}

group: ScienceData {

	group: Product {

	dimensions:
		mdrs                     = 30; // Nb of MDRs in this file
		nb_pixels                = UNLIMITED;
		time                     = 1;
		pixels_4_itime_1.5       = 4;
		pixels_4_itime_6         = 1;
		pixels_4_itime_0.1875    = 32;
		pixels_4_itime_0.0234375 = 256;
		corners                  = 4; // nb of corners
		// number of elements per bands
		rec_band_1A              = 659;  // seems to be fix for all band_1A recs if not they should be defined locally in each group
		rec_band_1B              = 365;  // same
		rec_band_2A              = 71;   // same
		rec_band_2B              = 953;  // same
		rec_band_3               = 1024; // same
		rec_band_4               = 1024; // same
		rec_band_5               = 15;   // same
		rec_band_6               = 15;   // same
		rec_band_shortPS         = 20;   // same
		rec_band_shortPP         = 20;   // same
		nb_itimes                = 6;    // max number of integration times
		unknown_dim = 3; // do not know why it is always 3

	variables:
		// in this case itimes will always be the max possible 6 and the number of pixels will be the max for all MDRs. The number of pixels used will determine which integration time had been used
		// the maximum integration time used for all MDRs in this file is for example 0.1875 which means that we need to have nb_pixels = 32 
		// Fill values are also going to be used a lot and the file size will be a little bit inflated but compression should be good.
		int start_time(mdrs,time) ;
			start_time:long_name = "reference time of a MDR" ;
			start_time:units     = "UTC time in epoch time: seconds since 1971 (epoc time)" ;

		int end_time(mdrs,time) ;
			end_time:long_name = "reference time of a MDR" ;
			end_time:units     = "UTC time in epoch time: seconds since 1971 (epoc time): seconds since 1971 (epoc time)" ;

		float itimes(mdrs, nb_itimes); // integration times
			itimes:long_name = "integration times";
			itimes:units     = "seconds" ;
			itimes:_FillValue = -999 ;
			itimes:valid_min = -127b ;
			itimes:valid_max = 127b ;

		float scanner_angle(mdrs, nb_itimes, pixels_4_itime_0.1875); // take the max of nb pixels for all possible integration times, need to use invalid values for not existing values
			scanner_angle:long_name  = "scanner angle";
			scanner_angle:units      = "degrees" ;
			scanner_angle:_FillValue = -999 ; 
			scanner_angle:valid_min  = -180 ; // QC values (example, not the right values)
			scanner_angle:valid_max  = 180  ; // QC values (example, not the right values)
	  
		float corners(mdrs, nb_itimes, corners, pixels_4_itime_0.1875); // take the max of nb pixels for all possible integration times, need to use invalid values for not existing values
			corners:long_name   = "pixel corners";
			corners:units       = "degrees";
			corners:_FillValue  = -999;
			corners:valid_min   = -180; // QC values (example, not the right values) 
			corners:valid_max   = 180; // QC values (example, not the right values) 

		float centers(mdrs, nb_itimes, pixels_4_itime_0.1875); // take the max of nb pixels for all possible integration times, need to use invalid values for not existing values (here it is 32 values)
			corners:long_name   = "pixel centre";
			corners:units       = "degrees";
			corners:_FillValue  = -999;
			corners:valid_min   = -180; // QC values (example, not the right values) 
			corners:valid_max   = 180; // QC values (example, not the right values) 

		float solar_zenith(mdrs, nb_itimes, unknown_dim, pixels_4_itime_0.1875); // same take the max possible number of pixels for all possible integration times (here 32 values)
			solar_zenith:long_name  = "solar zenith";
			solar_zenith:units      = "degrees";
			solar_zenith:_FillValue = -999;
			solar_zenith:valid_min  = -180; // QC values (example, not the right values) 
			solar_zenith:valid_max  = 180; // QC values (example, not the right values) 

		float wavelength_1A(mdrs, rec_band_1A);
			wavelength_1A:long_name  = "wavelength values for band 1A";
			wavelength_1A:units      = "nm";  
			wavelength_1A:_FillValue = -9999; // TBD
			wavelength_1A:valid_min  = 0; // TBD 
			wavelength_1A:valid_max  = 0; // TBD 

		float band_1A(mdrs, pixels_4_itime_0.1875, rec_band_1A); //a band is nb of pixels * nb of measures in a record
			band_1A:long_name  = "measures for band 1A";
			band_1A:units      = "BU";  // TBD
			band_1A:_FillValue = -9999; // TBD
			band_1A:valid_min  = 0; // TBD 
			band_1A:valid_max  = 0; // TBD 

		float wavelength_1B(mdrs, rec_band_1B);
			wavelength_1B:long_name  = "wavelength values for band 1B";
			wavelength_1B:units      = "nm";  
			wavelength_1B:_FillValue = -9999; // TBD
			wavelength_1B:valid_min  = 0; // TBD 
			wavelength_1A:valid_max  = 0; // TBD 

		float band_1B(mdrs, pixels_4_itime_0.1875,rec_band_1B); //a band is nb of pixels * nb of measures in a record
			band_1B:long_name  = "measures for band 1B";
			band_1B:units      = "BU";  // TBD
			band_1B:_FillValue = -9999; // TBD
			band_1B:valid_min  = 0; // TBD 
			band_1B:valid_max  = 0; // TBD 

		// Add the other bands
	  } // group Product
  } // Science Data

// global attributes:
 :Conventions = "CF-1.0" ;
 :title = "GOME ..." ;
 :DSD_entry_id = "" ;
 :references = "N/A" ;
 :institution = "EUMETSAT:copyright 2011 EUMETSAT" ;
 :contact = "Eumetsat help desk at http://www.eumetsat.int" ;
 :netcdf_version_id = "netcdf library version 4.1.1 of Dec  2 2010 14:09:08" ;
 :creation_date = "2011-04-29" ;
 :product_version = "0.2" ;
}
